module  module_name(
  input a,b,
  output x
);
endmodule
