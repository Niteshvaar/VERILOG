module or_g(
  input a,b,
  output x
);
  or o1(x,a,b);
endmodule
