module nor_g(
  input a,b,
  output x
);
  nor n1(x,a,b);
endmodule
