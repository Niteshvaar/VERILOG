module nand_g(
  input a,b,
  output x
);
  nand n1(x,a,b);
endmodule
