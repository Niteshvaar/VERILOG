module xnor_g(
  input a,b,
  output x
);
  xnor x1(x,a,b);
endmodule
