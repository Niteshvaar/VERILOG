module net_dec(
  input a,
  output x
);
  wire b;
  assign x=b;
endmodule
