module buffer(
  input a,
  output x
);
  buf b1(x,a);
endmodule
