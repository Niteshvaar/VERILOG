module not_g(
  input a,
  output x
);
  not n1(x,a);
endmodule
