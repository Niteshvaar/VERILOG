module and_g(
  input a,b,
  output x
);
  and a1(x,a,b);
endmodule
