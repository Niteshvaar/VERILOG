module xor_g(
  input a,b,
  output x
);
  xor x1(x,a,b);
endmodule
